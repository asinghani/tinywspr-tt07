/*
 * Copyright (c) 2024 Anish Singhani
 * SPDX-License-Identifier: Apache-2.0
 */

`default_nettype none

module tt_um_asinghani_tinywspr (
    input  wire [7:0] ui_in,    // Dedicated inputs
    output wire [7:0] uo_out,   // Dedicated outputs
    input  wire [7:0] uio_in,   // IOs: Input path
    output wire [7:0] uio_out,  // IOs: Output path
    output wire [7:0] uio_oe,   // IOs: Enable path (active high: 0=input, 1=output)
    input  wire       ena,      // always 1 when the design is powered, so you can ignore it
    input  wire       clk,      // clock
    input  wire       rst_n     // reset_n - low to reset
);

    assign uio_out = 0;
    assign uio_oe  = 0;

    reg config_start0, config_start1, config_start2;
    always @(posedge clk) begin
        config_start0 <= ui_in[1];
        config_start1 <= config_start0;
        config_start2 <= config_start1;
    end

    reg rf_start0, rf_start1, rf_start2;
    always @(posedge clk) begin
        rf_start0 <= ui_in[2];
        rf_start1 <= rf_start0;
        rf_start2 <= rf_start1;
    end

    reg config_valid0, config_valid1, config_valid2, config_validlast;
    always @(posedge clk) begin
        config_valid0 <= ui_in[0];
        config_valid1 <= config_valid0;
        config_valid2 <= config_valid1;
        config_validlast <= config_valid2;
    end

    TopLevel tl (
        .clock(clk),
        .reset(!rst_n),
        .io_config_bits_in(uio_in),
        .io_config_valid_in(config_valid2 && ~config_validlast),
        .io_config_start(config_start2),
        .io_rf_start(rf_start2),
        .io_rf_out(uo_out[0]),
        .io_bit_out(uo_out[7:6])
    )

    assign uo_out[1] = uo_out[0];
    assign uo_out[5:2] = 0;

endmodule
